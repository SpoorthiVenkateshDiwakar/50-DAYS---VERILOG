module tb;
