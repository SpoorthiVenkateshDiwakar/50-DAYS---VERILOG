module and_gate();
  input wire a,b;
  output reg y;
  assign y=a&b;
endmodule
