module half_adder;
